--+----------------------------------------------------------------------------
--|
--| NAMING CONVENSIONS :
--|
--|    xb_<port name>           = off-chip bidirectional port ( _pads file )
--|    xi_<port name>           = off-chip input port         ( _pads file )
--|    xo_<port name>           = off-chip output port        ( _pads file )
--|    b_<port name>            = on-chip bidirectional port
--|    i_<port name>            = on-chip input port
--|    o_<port name>            = on-chip output port
--|    c_<signal name>          = combinatorial signal
--|    f_<signal name>          = synchronous signal
--|    ff_<signal name>         = pipeline stage (ff_, fff_, etc.)
--|    <signal name>_n          = active low signal
--|    w_<signal name>          = top level wiring signal
--|    g_<generic name>         = generic
--|    k_<constant name>        = constant
--|    v_<variable name>        = variable
--|    sm_<state machine type>  = state machine type definition
--|    s_<signal name>          = state name
--|
--+----------------------------------------------------------------------------
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;


entity top_basys3 is
-- TODO
port(
        -- inputs
        clk     :   in std_logic; -- native 100MHz FPGA clock
        sw      :   in std_logic_vector(7 downto 0);
        btnU    :   in std_logic; -- master_reset
   --     btnL    :   in std_logic; -- clk_reset
     --   btnR    :   in std_logic; -- fsm_reset
        btnC    :   in std_logic; -- advance
        
        -- outputs
        led :   out std_logic_vector(15 downto 0);
        -- 7-segment display segments (active-low cathodes)
        seg :   out std_logic_vector(6 downto 0);
        -- 7-segment display active-low enables (anodes)
        an  :   out std_logic_vector(3 downto 0)
    );
end top_basys3;

architecture top_basys3_arch of top_basys3 is 
  
	-- declare components and signals
component sevenSegDecoder is
              port(
                 i_D : in std_logic_vector (3 downto 0);
                 o_S : out std_logic_vector (6 downto 0)--changed 7 from 6
              );    
            end component; 
            
component mux is
              port(
                 i_A : in std_logic_vector (7 downto 0);
                 i_B : in std_logic_vector (7 downto 0);
                 i_cycle : in std_logic_vector (3 downto 0);
                 i_result : in std_logic_vector (7 downto 0);
                 i_off : in std_logic_vector(7 downto 0); --set to ground, idk what this is tho
                 o_data : out std_logic_vector (7 downto 0)
              );    
            end component;            

component twoscomp_decimal is
              port(
                 i_binary : in std_logic_vector (7 downto 0);
                 o_negative : out std_logic_vector (3 downto 0);
                 o_hundreds : out std_logic_vector (3 downto 0);
                 o_tens : out std_logic_vector (3 downto 0);
                 o_ones : out std_logic_vector (3 downto 0)
              );    
            end component; 

component Controller_fsm is
              port(
                 i_adv : in std_logic;
                 i_reset : in std_logic;
                 i_clk : in std_logic;
                 o_cycle : out std_logic_vector (3 downto 0)
              );    
            end component; 

component reg is
              port(
                 i_operand : in std_logic_vector (7 downto 0);
                 i_fsm     : in std_logic_vector (3 downto 0);
                 o_operand : out std_logic_vector (7 downto 0)
              );    
            end component;             
            
component ALU is
              port(
                 i_A : in std_logic_vector (7 downto 0);
                 i_B : in std_logic_vector (7 downto 0);
                 i_op : in std_logic_vector (3 downto 0);
                 o_result : out std_logic_vector (7 downto 0);
                 o_carryOut : out std_logic_vector (2 downto 0)
              );    
            end component; 
                                       
component clock_divider is
            generic ( constant k_DIV : natural := 2    ); -- How many clk cycles until slow clock toggles
                                                       -- Effectively, you divide the clk double this 
                                                       -- number (e.g., k_DIV := 2 --> clock divider of 4)
            port (     i_clk    : in std_logic;
                    i_reset  : in std_logic;           -- asynchronous
                    o_clk    : out std_logic           -- divided (slow) clock
            );
        end component clock_divider;
                    
component TDM4 is
            generic ( constant k_WIDTH : natural  := 4); -- bits in input and output
            Port ( i_clk        : in  STD_LOGIC;
                   i_reset        : in  STD_LOGIC; -- asynchronous
                   i_D3         : in  STD_LOGIC_VECTOR (k_WIDTH - 1 downto 0);
                   i_D2         : in  STD_LOGIC_VECTOR (k_WIDTH - 1 downto 0);
                   i_D1         : in  STD_LOGIC_VECTOR (k_WIDTH - 1 downto 0);
                   i_D0         : in  STD_LOGIC_VECTOR (k_WIDTH - 1 downto 0);
                   o_data        : out STD_LOGIC_VECTOR (k_WIDTH - 1 downto 0);
                   o_sel        : out STD_LOGIC_VECTOR (3 downto 0)    -- selected data line (one-cold)
            );
        end component TDM4;
        
component regi is
            Port (
                    i_operand   : in std_logic_vector (7 downto 0);
                    i_cycle   : in std_logic_vector (3 downto 0);
                    o_operand   : out std_logic_vector (7 downto 0)
        );
        end component regi;
        
component regina is
            Port (
                    i_operand   : in std_logic_vector (7 downto 0);
                    i_cycle   : in std_logic_vector (3 downto 0);
                    o_operand   : out std_logic_vector (7 downto 0)
        );
                end component regina;
        --wires
        signal w_fsm : std_logic_vector(3 downto 0);
        signal w_clk : std_logic;
        signal w_A : std_logic_vector(7 downto 0);
        signal w_B : std_logic_vector(7 downto 0);
        signal w_ALU : std_logic_vector(7 downto 0);
        signal w_mux : std_logic_vector(7 downto 0);
        signal w_sign : std_logic_vector(3 downto 0);
        signal w_hund : std_logic_vector(3 downto 0);
        signal w_tens : std_logic_vector(3 downto 0);
        signal w_ones : std_logic_vector(3 downto 0);
        signal w_tdm : std_logic_vector(3 downto 0);
        signal w_btnU : std_logic;
        signal w_btnc : std_logic;
        
        --signals for registers?
        signal i_operand : std_logic_vector(7 downto 0);
        signal o_operand : std_logic_vector(7 downto 0);
        
        --signals for mux?
--        signal i_A : std_logic_vector(7 downto 0);
  --      signal i_B : std_logic_vector(7 downto 0);
    --    signal i_result : std_logic_vector(7 downto 0);
      --  signal i_cycle : std_logic_vector(7 downto 0);
       -- signal o_data : std_logic_vector(7 downto 0);
        
begin
	-- PORT MAPS ----------------------------------------
led(3 downto 0) <= w_fsm;
led(12 downto 4) <= "000000000";
w_btnU <= btnU;
w_btnC <= btnC;
	
regA_inst : regi port map (
                i_operand   => sw(7 downto 0),
                i_cycle     => w_fsm,
                o_operand   => w_A
    );
    
    regB_inst : regina port map (
                i_operand   => sw(7 downto 0),
                i_cycle     => w_fsm,
                o_operand   => w_B
    );


uut_inst : sevenSegDecoder port map (
               i_D     => w_tdm,
               o_S     => seg
           );
clkdiv_inst : clock_divider         --instantiation of clock_divider to take 
           generic map ( k_DIV => 50000000) -- 1 Hz clock from 100 MHz = 50mill
           port map (                          
               i_clk   => clk,
               i_reset => w_btnU,
               o_clk   => w_clk
           );  
	
tdm_inst : TDM4 --k_WIDTH needs help
          generic map ( k_WIDTH => 4) -- bits in input and output
          Port map ( i_clk  => w_clk,
             i_reset   => w_btnU, -- asynchronous
             i_D3      => w_sign,
             i_D2      => w_hund,
             i_D1      => w_tens,
             i_D0      => w_ones,
             o_data    => w_tdm,
             o_sel     => an   -- selected data line (one-cold)
              );
                  
controller_inst : Controller_fsm port map (
             i_reset     => w_btnU,
             i_adv       => w_btnC,
             i_clk       => clk,
             o_cycle     => w_fsm
                             );

ALU_inst : ALU port map (
             i_A       => w_A,
             i_B       => w_B,
             i_op      => sw(3 downto 0),
             o_result  => w_ALU,
             o_carryOut   => led(15 downto 13)  
              );     
twos_inst : twoscomp_decimal port map (
             i_binary       => w_mux,
             o_negative     => w_sign,
             o_hundreds     => w_hund,
             o_tens      => w_tens,
             o_ones      => w_ones
                );    


                                            
mux_inst : mux port map (
            i_A         => w_A,
            i_B         => w_B,
            i_result    => w_ALU,
            i_cycle     => w_fsm,
            o_data      => w_mux,
            i_off       => "00000000"
);        

                                    
	-- CONCURRENT STATEMENTS ----------------------------
	    --need to make mux in here but how??
	
	
-- PROCESSES --------------------------------------------------------------------
    -- state memory w/ asynchronous reset ---------------
    -----------------------------------------------------    
	
end top_basys3_arch;
